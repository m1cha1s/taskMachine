`timescale 1ns / 1ps

module lcdDriver(clk, e, data);

input clk;
output e;
output [2:0] data;



endmodule
