`timescale 1ns / 1ps

module interCoreCom(slowClk, medClk, fastClk);


endmodule
