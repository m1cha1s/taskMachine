`timescale 1ns / 1ps

module coreCommunicationController(fastClk, medClk);
input wire fastClk, medClk;

endmodule
